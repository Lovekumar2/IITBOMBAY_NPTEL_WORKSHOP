-- v_jtag.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity v_jtag is
	port (
		tck_clk                         : out std_logic;                                       --          tck.clk
		virtual_jtag_tdi                : out std_logic;                                       -- virtual_jtag.tdi
		virtual_jtag_tdo                : in  std_logic                    := '0';             --             .tdo
		virtual_jtag_ir_in              : out std_logic_vector(0 downto 0);                    --             .ir_in
		virtual_jtag_ir_out             : in  std_logic_vector(0 downto 0) := (others => '0'); --             .ir_out
		virtual_jtag_virtual_state_cdr  : out std_logic;                                       --             .virtual_state_cdr
		virtual_jtag_virtual_state_sdr  : out std_logic;                                       --             .virtual_state_sdr
		virtual_jtag_virtual_state_e1dr : out std_logic;                                       --             .virtual_state_e1dr
		virtual_jtag_virtual_state_pdr  : out std_logic;                                       --             .virtual_state_pdr
		virtual_jtag_virtual_state_e2dr : out std_logic;                                       --             .virtual_state_e2dr
		virtual_jtag_virtual_state_udr  : out std_logic;                                       --             .virtual_state_udr
		virtual_jtag_virtual_state_cir  : out std_logic;                                       --             .virtual_state_cir
		virtual_jtag_virtual_state_uir  : out std_logic;                                       --             .virtual_state_uir
		virtual_jtag_tms                : out std_logic;                                       --             .tms
		virtual_jtag_jtag_state_tlr     : out std_logic;                                       --             .jtag_state_tlr
		virtual_jtag_jtag_state_rti     : out std_logic;                                       --             .jtag_state_rti
		virtual_jtag_jtag_state_sdrs    : out std_logic;                                       --             .jtag_state_sdrs
		virtual_jtag_jtag_state_cdr     : out std_logic;                                       --             .jtag_state_cdr
		virtual_jtag_jtag_state_sdr     : out std_logic;                                       --             .jtag_state_sdr
		virtual_jtag_jtag_state_e1dr    : out std_logic;                                       --             .jtag_state_e1dr
		virtual_jtag_jtag_state_pdr     : out std_logic;                                       --             .jtag_state_pdr
		virtual_jtag_jtag_state_e2dr    : out std_logic;                                       --             .jtag_state_e2dr
		virtual_jtag_jtag_state_udr     : out std_logic;                                       --             .jtag_state_udr
		virtual_jtag_jtag_state_sirs    : out std_logic;                                       --             .jtag_state_sirs
		virtual_jtag_jtag_state_cir     : out std_logic;                                       --             .jtag_state_cir
		virtual_jtag_jtag_state_sir     : out std_logic;                                       --             .jtag_state_sir
		virtual_jtag_jtag_state_e1ir    : out std_logic;                                       --             .jtag_state_e1ir
		virtual_jtag_jtag_state_pir     : out std_logic;                                       --             .jtag_state_pir
		virtual_jtag_jtag_state_e2ir    : out std_logic;                                       --             .jtag_state_e2ir
		virtual_jtag_jtag_state_uir     : out std_logic                                        --             .jtag_state_uir
	);
end entity v_jtag;

architecture rtl of v_jtag is
	component sld_virtual_jtag is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			sld_ir_width            : integer := 1
		);
		port (
			tdi                : out std_logic;                                       -- tdi
			tdo                : in  std_logic                    := 'X';             -- tdo
			ir_in              : out std_logic_vector(0 downto 0);                    -- ir_in
			ir_out             : in  std_logic_vector(0 downto 0) := (others => 'X'); -- ir_out
			virtual_state_cdr  : out std_logic;                                       -- virtual_state_cdr
			virtual_state_sdr  : out std_logic;                                       -- virtual_state_sdr
			virtual_state_e1dr : out std_logic;                                       -- virtual_state_e1dr
			virtual_state_pdr  : out std_logic;                                       -- virtual_state_pdr
			virtual_state_e2dr : out std_logic;                                       -- virtual_state_e2dr
			virtual_state_udr  : out std_logic;                                       -- virtual_state_udr
			virtual_state_cir  : out std_logic;                                       -- virtual_state_cir
			virtual_state_uir  : out std_logic;                                       -- virtual_state_uir
			tms                : out std_logic;                                       -- tms
			jtag_state_tlr     : out std_logic;                                       -- jtag_state_tlr
			jtag_state_rti     : out std_logic;                                       -- jtag_state_rti
			jtag_state_sdrs    : out std_logic;                                       -- jtag_state_sdrs
			jtag_state_cdr     : out std_logic;                                       -- jtag_state_cdr
			jtag_state_sdr     : out std_logic;                                       -- jtag_state_sdr
			jtag_state_e1dr    : out std_logic;                                       -- jtag_state_e1dr
			jtag_state_pdr     : out std_logic;                                       -- jtag_state_pdr
			jtag_state_e2dr    : out std_logic;                                       -- jtag_state_e2dr
			jtag_state_udr     : out std_logic;                                       -- jtag_state_udr
			jtag_state_sirs    : out std_logic;                                       -- jtag_state_sirs
			jtag_state_cir     : out std_logic;                                       -- jtag_state_cir
			jtag_state_sir     : out std_logic;                                       -- jtag_state_sir
			jtag_state_e1ir    : out std_logic;                                       -- jtag_state_e1ir
			jtag_state_pir     : out std_logic;                                       -- jtag_state_pir
			jtag_state_e2ir    : out std_logic;                                       -- jtag_state_e2ir
			jtag_state_uir     : out std_logic;                                       -- jtag_state_uir
			tck                : out std_logic                                        -- clk
		);
	end component sld_virtual_jtag;

begin

	virtual_jtag_0 : component sld_virtual_jtag
		generic map (
			sld_auto_instance_index => "YES",
			sld_instance_index      => 0,
			sld_ir_width            => 1
		)
		port map (
			tdi                => virtual_jtag_tdi,                -- jtag.tdi
			tdo                => virtual_jtag_tdo,                --     .tdo
			ir_in              => virtual_jtag_ir_in,              --     .ir_in
			ir_out             => virtual_jtag_ir_out,             --     .ir_out
			virtual_state_cdr  => virtual_jtag_virtual_state_cdr,  --     .virtual_state_cdr
			virtual_state_sdr  => virtual_jtag_virtual_state_sdr,  --     .virtual_state_sdr
			virtual_state_e1dr => virtual_jtag_virtual_state_e1dr, --     .virtual_state_e1dr
			virtual_state_pdr  => virtual_jtag_virtual_state_pdr,  --     .virtual_state_pdr
			virtual_state_e2dr => virtual_jtag_virtual_state_e2dr, --     .virtual_state_e2dr
			virtual_state_udr  => virtual_jtag_virtual_state_udr,  --     .virtual_state_udr
			virtual_state_cir  => virtual_jtag_virtual_state_cir,  --     .virtual_state_cir
			virtual_state_uir  => virtual_jtag_virtual_state_uir,  --     .virtual_state_uir
			tms                => virtual_jtag_tms,                --     .tms
			jtag_state_tlr     => virtual_jtag_jtag_state_tlr,     --     .jtag_state_tlr
			jtag_state_rti     => virtual_jtag_jtag_state_rti,     --     .jtag_state_rti
			jtag_state_sdrs    => virtual_jtag_jtag_state_sdrs,    --     .jtag_state_sdrs
			jtag_state_cdr     => virtual_jtag_jtag_state_cdr,     --     .jtag_state_cdr
			jtag_state_sdr     => virtual_jtag_jtag_state_sdr,     --     .jtag_state_sdr
			jtag_state_e1dr    => virtual_jtag_jtag_state_e1dr,    --     .jtag_state_e1dr
			jtag_state_pdr     => virtual_jtag_jtag_state_pdr,     --     .jtag_state_pdr
			jtag_state_e2dr    => virtual_jtag_jtag_state_e2dr,    --     .jtag_state_e2dr
			jtag_state_udr     => virtual_jtag_jtag_state_udr,     --     .jtag_state_udr
			jtag_state_sirs    => virtual_jtag_jtag_state_sirs,    --     .jtag_state_sirs
			jtag_state_cir     => virtual_jtag_jtag_state_cir,     --     .jtag_state_cir
			jtag_state_sir     => virtual_jtag_jtag_state_sir,     --     .jtag_state_sir
			jtag_state_e1ir    => virtual_jtag_jtag_state_e1ir,    --     .jtag_state_e1ir
			jtag_state_pir     => virtual_jtag_jtag_state_pir,     --     .jtag_state_pir
			jtag_state_e2ir    => virtual_jtag_jtag_state_e2ir,    --     .jtag_state_e2ir
			jtag_state_uir     => virtual_jtag_jtag_state_uir,     --     .jtag_state_uir
			tck                => tck_clk                          --  tck.clk
		);

end architecture rtl; -- of v_jtag
